module RSstore(clock);
input clock;

always@(posedge clock)
begin
end

endmodule