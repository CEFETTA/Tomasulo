library verilog;
use verilog.vl_types.all;
entity RSload is
end RSload;
