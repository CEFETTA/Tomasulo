module RSadders(OP, Clock, Adderin, Busy);
  output reg Busy;
  reg [15:0] Qj, Qk, Vj, Vk;
  input [15:0] OP;
  input Clock, Adderin;
  
  
  
endmodule