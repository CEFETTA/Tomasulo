library verilog;
use verilog.vl_types.all;
entity RSstore is
end RSstore;
